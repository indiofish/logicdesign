`include "../alarm/AlarmModule.v"
`include "../stopwatch/StopWatch.v"
`include "../watch/Watch.v"
//add more extra implementation module's by include
`include "../stopwatch/SevenSegDecoder.v"

module WatchCtrl (

);
  
endmodule
