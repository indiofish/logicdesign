module D_flipflop(
  output Q, notQ,
  input D, CK
);

endmodule
